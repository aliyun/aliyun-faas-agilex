
`define Response_defaultEncoding_type [1:0]
`define Response_defaultEncoding_OKAY 2'b00
`define Response_defaultEncoding_RESERVED 2'b01
`define Response_defaultEncoding_SLAVEERROR 2'b10
`define Response_defaultEncoding_DECODEERROR 2'b11

