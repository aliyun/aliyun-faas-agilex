// ***************************************************************************************
//
// Filename        :    ddr_axi_cross_wrapper.v
// Projectname     :    F5
// Description     :                                             
// ***************************************************************************************
module  ddr4_axi4mm_cc_wrapper
#(
    parameter ADDR_WIDTH = 64 , 
    parameter DATA_WIDTH = 512,
    parameter WSTRB_WIDTH= 64  
)
(
    input                         kernel_clk            ,
    input                         kernel_clk_rst        ,

    input      [ADDR_WIDTH-1:0]   c0_sys_axi_araddr     ,
    input      [1:0]              c0_sys_axi_arburst    ,
    input      [3:0]              c0_sys_axi_arcache    ,
    input      [15:0]             c0_sys_axi_arid       ,
    input      [7:0]              c0_sys_axi_arlen      ,
    input      [0:0]              c0_sys_axi_arlock     ,
    input      [2:0]              c0_sys_axi_arprot     ,
    input      [3:0]              c0_sys_axi_arqos      ,
    output                        c0_sys_axi_arready    ,
    input      [3:0]              c0_sys_axi_arregion   ,
    input      [2:0]              c0_sys_axi_arsize     ,
    input                         c0_sys_axi_arvalid    ,
    input      [ADDR_WIDTH-1:0]   c0_sys_axi_awaddr     ,
    input      [1:0]              c0_sys_axi_awburst    ,
    input      [3:0]              c0_sys_axi_awcache    ,
    input      [15:0]             c0_sys_axi_awid       ,
    input      [7:0]              c0_sys_axi_awlen      ,
    input      [0:0]              c0_sys_axi_awlock     ,
    input      [2:0]              c0_sys_axi_awprot     ,
    input      [3:0]              c0_sys_axi_awqos      ,
    output                        c0_sys_axi_awready    ,
    input      [3:0]              c0_sys_axi_awregion   ,
    input      [2:0]              c0_sys_axi_awsize     ,
    input                         c0_sys_axi_awvalid    ,
    output     [15:0]             c0_sys_axi_bid        ,
    input                         c0_sys_axi_bready     ,
    output     [1:0]              c0_sys_axi_bresp      ,
    output                        c0_sys_axi_bvalid     ,
    output     [DATA_WIDTH-1:0]   c0_sys_axi_rdata      ,
    output     [15:0]             c0_sys_axi_rid        ,
    output                        c0_sys_axi_rlast      ,
    input                         c0_sys_axi_rready     ,
    output     [1:0]              c0_sys_axi_rresp      ,
    output                        c0_sys_axi_rvalid     ,
    input      [DATA_WIDTH-1:0]   c0_sys_axi_wdata      ,
    input                         c0_sys_axi_wlast      ,
    output                        c0_sys_axi_wready     ,
    input      [WSTRB_WIDTH-1:0]  c0_sys_axi_wstrb      ,
    input                         c0_sys_axi_wvalid     ,     

    input      [ADDR_WIDTH-1:0]   c1_sys_axi_araddr     ,
    input      [1:0]              c1_sys_axi_arburst    ,
    input      [3:0]              c1_sys_axi_arcache    ,
    input      [15:0]             c1_sys_axi_arid       ,
    input      [7:0]              c1_sys_axi_arlen      ,
    input      [0:0]              c1_sys_axi_arlock     ,
    input      [2:0]              c1_sys_axi_arprot     ,
    input      [3:0]              c1_sys_axi_arqos      ,
    output                        c1_sys_axi_arready    ,
    input      [3:0]              c1_sys_axi_arregion   ,
    input      [2:0]              c1_sys_axi_arsize     ,
    input                         c1_sys_axi_arvalid    ,
    input      [ADDR_WIDTH-1:0]   c1_sys_axi_awaddr     ,
    input      [1:0]              c1_sys_axi_awburst    ,
    input      [3:0]              c1_sys_axi_awcache    ,
    input      [15:0]             c1_sys_axi_awid       ,
    input      [7:0]              c1_sys_axi_awlen      ,
    input      [0:0]              c1_sys_axi_awlock     ,
    input      [2:0]              c1_sys_axi_awprot     ,
    input      [3:0]              c1_sys_axi_awqos      ,
    output                        c1_sys_axi_awready    ,
    input      [3:0]              c1_sys_axi_awregion   ,
    input      [2:0]              c1_sys_axi_awsize     ,
    input                         c1_sys_axi_awvalid    ,
    output     [15:0]             c1_sys_axi_bid        ,
    input                         c1_sys_axi_bready     ,
    output     [1:0]              c1_sys_axi_bresp      ,
    output                        c1_sys_axi_bvalid     ,
    output     [DATA_WIDTH-1:0]   c1_sys_axi_rdata      ,
    output     [15:0]             c1_sys_axi_rid        ,
    output                        c1_sys_axi_rlast      ,
    input                         c1_sys_axi_rready     ,
    output     [1:0]              c1_sys_axi_rresp      ,
    output                        c1_sys_axi_rvalid     ,
    input      [DATA_WIDTH-1:0]   c1_sys_axi_wdata      ,
    input                         c1_sys_axi_wlast      ,
    output                        c1_sys_axi_wready     ,
    input      [WSTRB_WIDTH-1:0]  c1_sys_axi_wstrb      ,
    input                         c1_sys_axi_wvalid     ,     

    input      [ADDR_WIDTH-1:0]   c2_sys_axi_araddr     ,
    input      [1:0]              c2_sys_axi_arburst    ,
    input      [3:0]              c2_sys_axi_arcache    ,
    input      [15:0]             c2_sys_axi_arid       ,
    input      [7:0]              c2_sys_axi_arlen      ,
    input      [0:0]              c2_sys_axi_arlock     ,
    input      [2:0]              c2_sys_axi_arprot     ,
    input      [3:0]              c2_sys_axi_arqos      ,
    output                        c2_sys_axi_arready    ,
    input      [3:0]              c2_sys_axi_arregion   ,
    input      [2:0]              c2_sys_axi_arsize     ,
    input                         c2_sys_axi_arvalid    ,
    input      [ADDR_WIDTH-1:0]   c2_sys_axi_awaddr     ,
    input      [1:0]              c2_sys_axi_awburst    ,
    input      [3:0]              c2_sys_axi_awcache    ,
    input      [15:0]             c2_sys_axi_awid       ,
    input      [7:0]              c2_sys_axi_awlen      ,
    input      [0:0]              c2_sys_axi_awlock     ,
    input      [2:0]              c2_sys_axi_awprot     ,
    input      [3:0]              c2_sys_axi_awqos      ,
    output                        c2_sys_axi_awready    ,
    input      [3:0]              c2_sys_axi_awregion   ,
    input      [2:0]              c2_sys_axi_awsize     ,
    input                         c2_sys_axi_awvalid    ,
    output     [15:0]             c2_sys_axi_bid        ,
    input                         c2_sys_axi_bready     ,
    output     [1:0]              c2_sys_axi_bresp      ,
    output                        c2_sys_axi_bvalid     ,
    output     [DATA_WIDTH-1:0]   c2_sys_axi_rdata      ,
    output     [15:0]             c2_sys_axi_rid        ,
    output                        c2_sys_axi_rlast      ,
    input                         c2_sys_axi_rready     ,
    output     [1:0]              c2_sys_axi_rresp      ,
    output                        c2_sys_axi_rvalid     ,
    input      [DATA_WIDTH-1:0]   c2_sys_axi_wdata      ,
    input                         c2_sys_axi_wlast      ,
    output                        c2_sys_axi_wready     ,
    input      [WSTRB_WIDTH-1:0]  c2_sys_axi_wstrb      ,
    input                         c2_sys_axi_wvalid     ,     

    input      [ADDR_WIDTH-1:0]   c3_sys_axi_araddr     ,
    input      [1:0]              c3_sys_axi_arburst    ,
    input      [3:0]              c3_sys_axi_arcache    ,
    input      [15:0]             c3_sys_axi_arid       ,
    input      [7:0]              c3_sys_axi_arlen      ,
    input      [0:0]              c3_sys_axi_arlock     ,
    input      [2:0]              c3_sys_axi_arprot     ,
    input      [3:0]              c3_sys_axi_arqos      ,
    output                        c3_sys_axi_arready    ,
    input      [3:0]              c3_sys_axi_arregion   ,
    input      [2:0]              c3_sys_axi_arsize     ,
    input                         c3_sys_axi_arvalid    ,
    input      [ADDR_WIDTH-1:0]   c3_sys_axi_awaddr     ,
    input      [1:0]              c3_sys_axi_awburst    ,
    input      [3:0]              c3_sys_axi_awcache    ,
    input      [15:0]             c3_sys_axi_awid       ,
    input      [7:0]              c3_sys_axi_awlen      ,
    input      [0:0]              c3_sys_axi_awlock     ,
    input      [2:0]              c3_sys_axi_awprot     ,
    input      [3:0]              c3_sys_axi_awqos      ,
    output                        c3_sys_axi_awready    ,
    input      [3:0]              c3_sys_axi_awregion   ,
    input      [2:0]              c3_sys_axi_awsize     ,
    input                         c3_sys_axi_awvalid    ,
    output     [15:0]             c3_sys_axi_bid        ,
    input                         c3_sys_axi_bready     ,
    output     [1:0]              c3_sys_axi_bresp      ,
    output                        c3_sys_axi_bvalid     ,
    output     [DATA_WIDTH-1:0]   c3_sys_axi_rdata      ,
    output     [15:0]             c3_sys_axi_rid        ,
    output                        c3_sys_axi_rlast      ,
    input                         c3_sys_axi_rready     ,
    output     [1:0]              c3_sys_axi_rresp      ,
    output                        c3_sys_axi_rvalid     ,
    input      [DATA_WIDTH-1:0]   c3_sys_axi_wdata      ,
    input                         c3_sys_axi_wlast      ,
    output                        c3_sys_axi_wready     ,
    input      [WSTRB_WIDTH-1:0]  c3_sys_axi_wstrb      ,
    input                         c3_sys_axi_wvalid     ,     
 
    input                         c0_ddr4_usr_reset       ,   
    input                         c0_ddr4_usr_clk         ,   
    output     [63:0]             c0_ddr4_axi_araddr      ,
    output     [1:0]              c0_ddr4_axi_arburst     ,
    output     [3:0]              c0_ddr4_axi_arcache     ,
    output     [4:0]              c0_ddr4_axi_arid        ,
    output     [7:0]              c0_ddr4_axi_arlen       ,
    output     [0:0]              c0_ddr4_axi_arlock      ,
    output     [2:0]              c0_ddr4_axi_arprot      ,
    output     [3:0]              c0_ddr4_axi_arqos       ,
    input                         c0_ddr4_axi_arready     ,
    output     [3:0]              c0_ddr4_axi_arregion    ,
    output     [2:0]              c0_ddr4_axi_arsize      ,
    output                        c0_ddr4_axi_arvalid     ,
    output     [63:0]             c0_ddr4_axi_awaddr      ,
    output     [1:0]              c0_ddr4_axi_awburst     ,
    output     [3:0]              c0_ddr4_axi_awcache     ,
    output     [4:0]              c0_ddr4_axi_awid        ,
    output     [7:0]              c0_ddr4_axi_awlen       ,
    output     [0:0]              c0_ddr4_axi_awlock      ,
    output     [2:0]              c0_ddr4_axi_awprot      ,
    output     [3:0]              c0_ddr4_axi_awqos       ,
    input                         c0_ddr4_axi_awready     ,
    output     [3:0]              c0_ddr4_axi_awregion    ,
    output     [2:0]              c0_ddr4_axi_awsize      ,
    output                        c0_ddr4_axi_awvalid     ,
    input      [4:0]              c0_ddr4_axi_bid         ,
    output                        c0_ddr4_axi_bready      ,
    input      [1:0]              c0_ddr4_axi_bresp       ,
    input                         c0_ddr4_axi_bvalid      ,
    input      [511:0]            c0_ddr4_axi_rdata       ,
    input      [4:0]              c0_ddr4_axi_rid         ,
    input                         c0_ddr4_axi_rlast       ,
    output                        c0_ddr4_axi_rready      ,
    input      [1:0]              c0_ddr4_axi_rresp       ,
    input                         c0_ddr4_axi_rvalid      ,
    output     [511:0]            c0_ddr4_axi_wdata       ,
    output                        c0_ddr4_axi_wlast       ,
    input                         c0_ddr4_axi_wready      ,
    output     [63:0]             c0_ddr4_axi_wstrb       ,
    output                        c0_ddr4_axi_wvalid      ,     
    
    input                         c1_ddr4_usr_reset      ,   
    input                         c1_ddr4_usr_clk        ,   
    output     [63:0]             c1_ddr4_axi_araddr      ,
    output     [1:0]              c1_ddr4_axi_arburst     ,
    output     [3:0]              c1_ddr4_axi_arcache     ,
    output     [4:0]              c1_ddr4_axi_arid        ,
    output     [7:0]              c1_ddr4_axi_arlen       ,
    output     [0:0]              c1_ddr4_axi_arlock      ,
    output     [2:0]              c1_ddr4_axi_arprot      ,
    output     [3:0]              c1_ddr4_axi_arqos       ,
    input                         c1_ddr4_axi_arready     ,
    output     [3:0]              c1_ddr4_axi_arregion    ,
    output     [2:0]              c1_ddr4_axi_arsize      ,
    output                        c1_ddr4_axi_arvalid     ,
    output     [63:0]             c1_ddr4_axi_awaddr      ,
    output     [1:0]              c1_ddr4_axi_awburst     ,
    output     [3:0]              c1_ddr4_axi_awcache     ,
    output     [4:0]              c1_ddr4_axi_awid        ,
    output     [7:0]              c1_ddr4_axi_awlen       ,
    output     [0:0]              c1_ddr4_axi_awlock      ,
    output     [2:0]              c1_ddr4_axi_awprot      ,
    output     [3:0]              c1_ddr4_axi_awqos       ,
    input                         c1_ddr4_axi_awready     ,
    output     [3:0]              c1_ddr4_axi_awregion    ,
    output     [2:0]              c1_ddr4_axi_awsize      ,
    output                        c1_ddr4_axi_awvalid     ,
    input      [4:0]              c1_ddr4_axi_bid         ,
    output                        c1_ddr4_axi_bready      ,
    input      [1:0]              c1_ddr4_axi_bresp       ,
    input                         c1_ddr4_axi_bvalid      ,
    input      [511:0]            c1_ddr4_axi_rdata       ,
    input      [4:0]              c1_ddr4_axi_rid         ,
    input                         c1_ddr4_axi_rlast       ,
    output                        c1_ddr4_axi_rready      ,
    input      [1:0]              c1_ddr4_axi_rresp       ,
    input                         c1_ddr4_axi_rvalid      ,
    output     [511:0]            c1_ddr4_axi_wdata       ,
    output                        c1_ddr4_axi_wlast       ,
    input                         c1_ddr4_axi_wready      ,
    output     [63:0]             c1_ddr4_axi_wstrb       ,
    output                        c1_ddr4_axi_wvalid      ,

    input                         c2_ddr4_usr_reset       ,   
    input                         c2_ddr4_usr_clk         ,   
    output     [63:0]             c2_ddr4_axi_araddr      ,
    output     [1:0]              c2_ddr4_axi_arburst     ,
    output     [3:0]              c2_ddr4_axi_arcache     ,
    output     [4:0]              c2_ddr4_axi_arid        ,
    output     [7:0]              c2_ddr4_axi_arlen       ,
    output     [0:0]              c2_ddr4_axi_arlock      ,
    output     [2:0]              c2_ddr4_axi_arprot      ,
    output     [3:0]              c2_ddr4_axi_arqos       ,
    input                         c2_ddr4_axi_arready     ,
    output     [3:0]              c2_ddr4_axi_arregion    ,
    output     [2:0]              c2_ddr4_axi_arsize      ,
    output                        c2_ddr4_axi_arvalid     ,
    output     [63:0]             c2_ddr4_axi_awaddr      ,
    output     [1:0]              c2_ddr4_axi_awburst     ,
    output     [3:0]              c2_ddr4_axi_awcache     ,
    output     [4:0]              c2_ddr4_axi_awid        ,
    output     [7:0]              c2_ddr4_axi_awlen       ,
    output     [0:0]              c2_ddr4_axi_awlock      ,
    output     [2:0]              c2_ddr4_axi_awprot      ,
    output     [3:0]              c2_ddr4_axi_awqos       ,
    input                         c2_ddr4_axi_awready     ,
    output     [3:0]              c2_ddr4_axi_awregion    ,
    output     [2:0]              c2_ddr4_axi_awsize      ,
    output                        c2_ddr4_axi_awvalid     ,
    input      [4:0]              c2_ddr4_axi_bid         ,
    output                        c2_ddr4_axi_bready      ,
    input      [1:0]              c2_ddr4_axi_bresp       ,
    input                         c2_ddr4_axi_bvalid      ,
    input      [511:0]            c2_ddr4_axi_rdata       ,
    input      [4:0]              c2_ddr4_axi_rid         ,
    input                         c2_ddr4_axi_rlast       ,
    output                        c2_ddr4_axi_rready      ,
    input      [1:0]              c2_ddr4_axi_rresp       ,
    input                         c2_ddr4_axi_rvalid      ,
    output     [511:0]            c2_ddr4_axi_wdata       ,
    output                        c2_ddr4_axi_wlast       ,
    input                         c2_ddr4_axi_wready      ,
    output     [63:0]             c2_ddr4_axi_wstrb       ,
    output                        c2_ddr4_axi_wvalid      ,

    input                         c3_ddr4_usr_reset       ,   
    input                         c3_ddr4_usr_clk         ,   
    output     [63:0]             c3_ddr4_axi_araddr      ,
    output     [1:0]              c3_ddr4_axi_arburst     ,
    output     [3:0]              c3_ddr4_axi_arcache     ,
    output     [4:0]              c3_ddr4_axi_arid        ,
    output     [7:0]              c3_ddr4_axi_arlen       ,
    output     [0:0]              c3_ddr4_axi_arlock      ,
    output     [2:0]              c3_ddr4_axi_arprot      ,
    output     [3:0]              c3_ddr4_axi_arqos       ,
    input                         c3_ddr4_axi_arready     ,
    output     [3:0]              c3_ddr4_axi_arregion    ,
    output     [2:0]              c3_ddr4_axi_arsize      ,
    output                        c3_ddr4_axi_arvalid     ,
    output     [63:0]             c3_ddr4_axi_awaddr      ,
    output     [1:0]              c3_ddr4_axi_awburst     ,
    output     [3:0]              c3_ddr4_axi_awcache     ,
    output     [4:0]              c3_ddr4_axi_awid        ,
    output     [7:0]              c3_ddr4_axi_awlen       ,
    output     [0:0]              c3_ddr4_axi_awlock      ,
    output     [2:0]              c3_ddr4_axi_awprot      ,
    output     [3:0]              c3_ddr4_axi_awqos       ,
    input                         c3_ddr4_axi_awready     ,
    output     [3:0]              c3_ddr4_axi_awregion    ,
    output     [2:0]              c3_ddr4_axi_awsize      ,
    output                        c3_ddr4_axi_awvalid     ,
    input      [4:0]              c3_ddr4_axi_bid         ,
    output                        c3_ddr4_axi_bready      ,
    input      [1:0]              c3_ddr4_axi_bresp       ,
    input                         c3_ddr4_axi_bvalid      ,
    input      [511:0]            c3_ddr4_axi_rdata       ,
    input      [4:0]              c3_ddr4_axi_rid         ,
    input                         c3_ddr4_axi_rlast       ,
    output                        c3_ddr4_axi_rready      ,
    input      [1:0]              c3_ddr4_axi_rresp       ,
    input                         c3_ddr4_axi_rvalid      ,
    output     [511:0]            c3_ddr4_axi_wdata       ,
    output                        c3_ddr4_axi_wlast       ,
    input                         c3_ddr4_axi_wready      ,
    output     [63:0]             c3_ddr4_axi_wstrb       ,
    output                        c3_ddr4_axi_wvalid
);

// ---------------------------------------------------------------------------------------
//  parameter
// ---------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------
//  signales
// ---------------------------------------------------------------------------------------

// ---------------------------------------------------------------------------------------
//  logic
// ---------------------------------------------------------------------------------------
ddr4_mmAxi4CC_std     c0_Axi4CCByToggle 
(
    .input_awvalid    (c0_sys_axi_awvalid  ),
    .input_awready    (c0_sys_axi_awready  ),
    .input_awaddr     (c0_sys_axi_awaddr   ),
    .input_awid       (c0_sys_axi_awid     ),
    .input_awlen      (c0_sys_axi_awlen    ),
    .input_awsize     (c0_sys_axi_awsize   ),
    .input_awburst    (c0_sys_axi_awburst  ),
    .input_wvalid     (c0_sys_axi_wvalid   ),
    .input_wready     (c0_sys_axi_wready   ),
    .input_wdata      (c0_sys_axi_wdata    ),
    .input_wstrb      (c0_sys_axi_wstrb    ),
    .input_wlast      (c0_sys_axi_wlast    ),
    .input_bvalid     (c0_sys_axi_bvalid   ),
    .input_bready     (c0_sys_axi_bready   ),
    .input_bid        (c0_sys_axi_bid      ),
    .input_bresp      (c0_sys_axi_bresp    ),
    .input_arvalid    (c0_sys_axi_arvalid  ),
    .input_arready    (c0_sys_axi_arready  ),
    .input_araddr     (c0_sys_axi_araddr   ),
    .input_arid       (c0_sys_axi_arid     ),
    .input_arlen      (c0_sys_axi_arlen    ),
    .input_arsize     (c0_sys_axi_arsize   ),
    .input_arburst    (c0_sys_axi_arburst  ),
    .input_rvalid     (c0_sys_axi_rvalid   ),
    .input_rready     (c0_sys_axi_rready   ),
    .input_rdata      (c0_sys_axi_rdata    ),
    .input_rid        (c0_sys_axi_rid      ),
    .input_rresp      (c0_sys_axi_rresp    ),
    .input_rlast      (c0_sys_axi_rlast    ),
    .output_awvalid   (c0_ddr4_axi_awvalid ),
    .output_awready   (c0_ddr4_axi_awready ),
    .output_awaddr    (c0_ddr4_axi_awaddr  ),
    .output_awid      (c0_ddr4_axi_awid    ),
    .output_awlen     (c0_ddr4_axi_awlen   ),
    .output_awsize    (c0_ddr4_axi_awsize  ),
    .output_awburst   (c0_ddr4_axi_awburst ),
    .output_wvalid    (c0_ddr4_axi_wvalid  ),
    .output_wready    (c0_ddr4_axi_wready  ),
    .output_wdata     (c0_ddr4_axi_wdata   ),
    .output_wstrb     (c0_ddr4_axi_wstrb   ),
    .output_wlast     (c0_ddr4_axi_wlast   ),
    .output_bvalid    (c0_ddr4_axi_bvalid  ),
    .output_bready    (c0_ddr4_axi_bready  ),
    .output_bid       (c0_ddr4_axi_bid     ),
    .output_bresp     (c0_ddr4_axi_bresp   ),
    .output_arvalid   (c0_ddr4_axi_arvalid ),
    .output_arready   (c0_ddr4_axi_arready ),
    .output_araddr    (c0_ddr4_axi_araddr  ),
    .output_arid      (c0_ddr4_axi_arid    ),
    .output_arlen     (c0_ddr4_axi_arlen   ),
    .output_arsize    (c0_ddr4_axi_arsize  ),
    .output_arburst   (c0_ddr4_axi_arburst ),
    .output_rvalid    (c0_ddr4_axi_rvalid  ),
    .output_rready    (c0_ddr4_axi_rready  ),
    .output_rdata     (c0_ddr4_axi_rdata   ),
    .output_rid       (c0_ddr4_axi_rid     ),
    .output_rresp     (c0_ddr4_axi_rresp   ),
    .output_rlast     (c0_ddr4_axi_rlast   ),
    .clkA_clk         (kernel_clk          ),
    .clkA_reset       (kernel_clk_rst      ),
    .clkB_clk         (c0_ddr4_usr_clk     ),
    .clkB_reset       (c0_ddr4_usr_reset   )
);

ddr4_mmAxi4CC_std    c1_Axi4CCByToggle 
(
    .input_awvalid    (c1_sys_axi_awvalid  ),
    .input_awready    (c1_sys_axi_awready  ),
    .input_awaddr     (c1_sys_axi_awaddr   ),
    .input_awid       (c1_sys_axi_awid     ),
    .input_awlen      (c1_sys_axi_awlen    ),
    .input_awsize     (c1_sys_axi_awsize   ),
    .input_awburst    (c1_sys_axi_awburst  ),
    .input_wvalid     (c1_sys_axi_wvalid   ),
    .input_wready     (c1_sys_axi_wready   ),
    .input_wdata      (c1_sys_axi_wdata    ),
    .input_wstrb      (c1_sys_axi_wstrb    ),
    .input_wlast      (c1_sys_axi_wlast    ),
    .input_bvalid     (c1_sys_axi_bvalid   ),
    .input_bready     (c1_sys_axi_bready   ),
    .input_bid        (c1_sys_axi_bid      ),
    .input_bresp      (c1_sys_axi_bresp    ),
    .input_arvalid    (c1_sys_axi_arvalid  ),
    .input_arready    (c1_sys_axi_arready  ),
    .input_araddr     (c1_sys_axi_araddr   ),
    .input_arid       (c1_sys_axi_arid     ),
    .input_arlen      (c1_sys_axi_arlen    ),
    .input_arsize     (c1_sys_axi_arsize   ),
    .input_arburst    (c1_sys_axi_arburst  ),
    .input_rvalid     (c1_sys_axi_rvalid   ),
    .input_rready     (c1_sys_axi_rready   ),
    .input_rdata      (c1_sys_axi_rdata    ),
    .input_rid        (c1_sys_axi_rid      ),
    .input_rresp      (c1_sys_axi_rresp    ),
    .input_rlast      (c1_sys_axi_rlast    ),
    .output_awvalid   (c1_ddr4_axi_awvalid ),
    .output_awready   (c1_ddr4_axi_awready ),
    .output_awaddr    (c1_ddr4_axi_awaddr  ),
    .output_awid      (c1_ddr4_axi_awid    ),
    .output_awlen     (c1_ddr4_axi_awlen   ),
    .output_awsize    (c1_ddr4_axi_awsize  ),
    .output_awburst   (c1_ddr4_axi_awburst ),
    .output_wvalid    (c1_ddr4_axi_wvalid  ),
    .output_wready    (c1_ddr4_axi_wready  ),
    .output_wdata     (c1_ddr4_axi_wdata   ),
    .output_wstrb     (c1_ddr4_axi_wstrb   ),
    .output_wlast     (c1_ddr4_axi_wlast   ),
    .output_bvalid    (c1_ddr4_axi_bvalid  ),
    .output_bready    (c1_ddr4_axi_bready  ),
    .output_bid       (c1_ddr4_axi_bid     ),
    .output_bresp     (c1_ddr4_axi_bresp   ),
    .output_arvalid   (c1_ddr4_axi_arvalid ),
    .output_arready   (c1_ddr4_axi_arready ),
    .output_araddr    (c1_ddr4_axi_araddr  ),
    .output_arid      (c1_ddr4_axi_arid    ),
    .output_arlen     (c1_ddr4_axi_arlen   ),
    .output_arsize    (c1_ddr4_axi_arsize  ),
    .output_arburst   (c1_ddr4_axi_arburst ),
    .output_rvalid    (c1_ddr4_axi_rvalid  ),
    .output_rready    (c1_ddr4_axi_rready  ),
    .output_rdata     (c1_ddr4_axi_rdata   ),
    .output_rid       (c1_ddr4_axi_rid     ),
    .output_rresp     (c1_ddr4_axi_rresp   ),
    .output_rlast     (c1_ddr4_axi_rlast   ),
    .clkA_clk         (kernel_clk          ),
    .clkA_reset       (kernel_clk_rst      ),
    .clkB_clk         (c1_ddr4_usr_clk     ),
    .clkB_reset       (c1_ddr4_usr_reset  )
);

ddr4_mmAxi4CC_std    c2_Axi4CCByToggle 
(
    .input_awvalid    (c2_sys_axi_awvalid  ),
    .input_awready    (c2_sys_axi_awready  ),
    .input_awaddr     (c2_sys_axi_awaddr   ),
    .input_awid       (c2_sys_axi_awid     ),
    .input_awlen      (c2_sys_axi_awlen    ),
    .input_awsize     (c2_sys_axi_awsize   ),
    .input_awburst    (c2_sys_axi_awburst  ),
    .input_wvalid     (c2_sys_axi_wvalid   ),
    .input_wready     (c2_sys_axi_wready   ),
    .input_wdata      (c2_sys_axi_wdata    ),
    .input_wstrb      (c2_sys_axi_wstrb    ),
    .input_wlast      (c2_sys_axi_wlast    ),
    .input_bvalid     (c2_sys_axi_bvalid   ),
    .input_bready     (c2_sys_axi_bready   ),
    .input_bid        (c2_sys_axi_bid      ),
    .input_bresp      (c2_sys_axi_bresp    ),
    .input_arvalid    (c2_sys_axi_arvalid  ),
    .input_arready    (c2_sys_axi_arready  ),
    .input_araddr     (c2_sys_axi_araddr   ),
    .input_arid       (c2_sys_axi_arid     ),
    .input_arlen      (c2_sys_axi_arlen    ),
    .input_arsize     (c2_sys_axi_arsize   ),
    .input_arburst    (c2_sys_axi_arburst  ),
    .input_rvalid     (c2_sys_axi_rvalid   ),
    .input_rready     (c2_sys_axi_rready   ),
    .input_rdata      (c2_sys_axi_rdata    ),
    .input_rid        (c2_sys_axi_rid      ),
    .input_rresp      (c2_sys_axi_rresp    ),
    .input_rlast      (c2_sys_axi_rlast    ),
    .output_awvalid   (c2_ddr4_axi_awvalid ),
    .output_awready   (c2_ddr4_axi_awready ),
    .output_awaddr    (c2_ddr4_axi_awaddr  ),
    .output_awid      (c2_ddr4_axi_awid    ),
    .output_awlen     (c2_ddr4_axi_awlen   ),
    .output_awsize    (c2_ddr4_axi_awsize  ),
    .output_awburst   (c2_ddr4_axi_awburst ),
    .output_wvalid    (c2_ddr4_axi_wvalid  ),
    .output_wready    (c2_ddr4_axi_wready  ),
    .output_wdata     (c2_ddr4_axi_wdata   ),
    .output_wstrb     (c2_ddr4_axi_wstrb   ),
    .output_wlast     (c2_ddr4_axi_wlast   ),
    .output_bvalid    (c2_ddr4_axi_bvalid  ),
    .output_bready    (c2_ddr4_axi_bready  ),
    .output_bid       (c2_ddr4_axi_bid     ),
    .output_bresp     (c2_ddr4_axi_bresp   ),
    .output_arvalid   (c2_ddr4_axi_arvalid ),
    .output_arready   (c2_ddr4_axi_arready ),
    .output_araddr    (c2_ddr4_axi_araddr  ),
    .output_arid      (c2_ddr4_axi_arid    ),
    .output_arlen     (c2_ddr4_axi_arlen   ),
    .output_arsize    (c2_ddr4_axi_arsize  ),
    .output_arburst   (c2_ddr4_axi_arburst ),
    .output_rvalid    (c2_ddr4_axi_rvalid  ),
    .output_rready    (c2_ddr4_axi_rready  ),
    .output_rdata     (c2_ddr4_axi_rdata   ),
    .output_rid       (c2_ddr4_axi_rid     ),
    .output_rresp     (c2_ddr4_axi_rresp   ),
    .output_rlast     (c2_ddr4_axi_rlast   ),
    .clkA_clk         (kernel_clk          ),
    .clkA_reset       (kernel_clk_rst      ),
    .clkB_clk         (c2_ddr4_usr_clk     ),
    .clkB_reset       (c2_ddr4_usr_reset   )
);

ddr4_mmAxi4CC_std     c3_Axi4CCByToggle 
(
    .input_awvalid    (c3_sys_axi_awvalid  ),
    .input_awready    (c3_sys_axi_awready  ),
    .input_awaddr     (c3_sys_axi_awaddr   ),
    .input_awid       (c3_sys_axi_awid     ),
    .input_awlen      (c3_sys_axi_awlen    ),
    .input_awsize     (c3_sys_axi_awsize   ),
    .input_awburst    (c3_sys_axi_awburst  ),
    .input_wvalid     (c3_sys_axi_wvalid   ),
    .input_wready     (c3_sys_axi_wready   ),
    .input_wdata      (c3_sys_axi_wdata    ),
    .input_wstrb      (c3_sys_axi_wstrb    ),
    .input_wlast      (c3_sys_axi_wlast    ),
    .input_bvalid     (c3_sys_axi_bvalid   ),
    .input_bready     (c3_sys_axi_bready   ),
    .input_bid        (c3_sys_axi_bid      ),
    .input_bresp      (c3_sys_axi_bresp    ),
    .input_arvalid    (c3_sys_axi_arvalid  ),
    .input_arready    (c3_sys_axi_arready  ),
    .input_araddr     (c3_sys_axi_araddr   ),
    .input_arid       (c3_sys_axi_arid     ),
    .input_arlen      (c3_sys_axi_arlen    ),
    .input_arsize     (c3_sys_axi_arsize   ),
    .input_arburst    (c3_sys_axi_arburst  ),
    .input_rvalid     (c3_sys_axi_rvalid   ),
    .input_rready     (c3_sys_axi_rready   ),
    .input_rdata      (c3_sys_axi_rdata    ),
    .input_rid        (c3_sys_axi_rid      ),
    .input_rresp      (c3_sys_axi_rresp    ),
    .input_rlast      (c3_sys_axi_rlast    ),
    .output_awvalid   (c3_ddr4_axi_awvalid ),
    .output_awready   (c3_ddr4_axi_awready ),
    .output_awaddr    (c3_ddr4_axi_awaddr  ),
    .output_awid      (c3_ddr4_axi_awid    ),
    .output_awlen     (c3_ddr4_axi_awlen   ),
    .output_awsize    (c3_ddr4_axi_awsize  ),
    .output_awburst   (c3_ddr4_axi_awburst ),
    .output_wvalid    (c3_ddr4_axi_wvalid  ),
    .output_wready    (c3_ddr4_axi_wready  ),
    .output_wdata     (c3_ddr4_axi_wdata   ),
    .output_wstrb     (c3_ddr4_axi_wstrb   ),
    .output_wlast     (c3_ddr4_axi_wlast   ),
    .output_bvalid    (c3_ddr4_axi_bvalid  ),
    .output_bready    (c3_ddr4_axi_bready  ),
    .output_bid       (c3_ddr4_axi_bid     ),
    .output_bresp     (c3_ddr4_axi_bresp   ),
    .output_arvalid   (c3_ddr4_axi_arvalid ),
    .output_arready   (c3_ddr4_axi_arready ),
    .output_araddr    (c3_ddr4_axi_araddr  ),
    .output_arid      (c3_ddr4_axi_arid    ),
    .output_arlen     (c3_ddr4_axi_arlen   ),
    .output_arsize    (c3_ddr4_axi_arsize  ),
    .output_arburst   (c3_ddr4_axi_arburst ),
    .output_rvalid    (c3_ddr4_axi_rvalid  ),
    .output_rready    (c3_ddr4_axi_rready  ),
    .output_rdata     (c3_ddr4_axi_rdata   ),
    .output_rid       (c3_ddr4_axi_rid     ),
    .output_rresp     (c3_ddr4_axi_rresp   ),
    .output_rlast     (c3_ddr4_axi_rlast   ),
    .clkA_clk         (kernel_clk          ),
    .clkA_reset       (kernel_clk_rst      ),
    .clkB_clk         (c3_ddr4_usr_clk     ),
    .clkB_reset       (c3_ddr4_usr_reset   )
);

endmodule
